package ram_constants is
	constant DATA_WIDTH : integer := 256;
	constant ADDR_WIDTH : integer := 8;
end package ram_constants;